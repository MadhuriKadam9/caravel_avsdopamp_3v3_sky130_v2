magic
tech sky130A
timestamp 1633972554
<< nwell >>
rect -1550 784 1272 1490
rect -1541 -1027 1263 784
<< pmos >>
rect -1293 -160 996 107
<< pdiff >>
rect -1293 565 996 708
rect -1293 308 -1083 565
rect -816 555 996 565
rect -816 308 490 555
rect -1293 298 490 308
rect 757 298 996 555
rect -1293 107 996 298
rect -1293 -341 996 -160
rect -1293 -370 500 -341
rect -1293 -627 -1083 -370
rect -816 -598 500 -370
rect 767 -598 996 -341
rect -816 -627 996 -598
rect -1293 -703 996 -627
<< pdiffc >>
rect -1083 308 -816 565
rect 490 298 757 555
rect -1083 -627 -816 -370
rect 500 -598 767 -341
<< nsubdiff >>
rect -1312 1109 1005 1242
rect -1312 880 -1073 1109
rect -816 880 1005 1109
rect -1312 737 1005 880
<< nsubdiffcont >>
rect -1073 880 -816 1109
<< poly >>
rect -1779 -160 -1293 107
rect 996 -160 1606 107
<< locali >>
rect -1321 1109 996 1242
rect -1321 1106 -1073 1109
rect -1321 879 -1076 1106
rect -816 880 996 1109
rect -819 879 996 880
rect -1321 565 996 879
rect -1321 556 -1083 565
rect -1312 308 -1083 556
rect -816 555 996 565
rect -816 308 490 555
rect -1312 298 490 308
rect 757 298 996 555
rect -1312 174 996 298
rect -1312 -341 996 -226
rect -1312 -370 500 -341
rect -1312 -627 -1083 -370
rect -816 -598 500 -370
rect 767 -598 996 -341
rect -816 -627 996 -598
rect -1312 -703 996 -627
<< viali >>
rect -1076 880 -1073 1106
rect -1073 880 -819 1106
rect -1076 879 -819 880
<< metal1 >>
rect -1317 1106 998 1249
rect -1317 879 -1076 1106
rect -819 879 998 1106
rect -1317 729 998 879
<< end >>
