magic
tech sky130A
timestamp 1634047645
<< nwell >>
rect 5589 5668 6996 6290
rect 11240 5731 12532 6097
rect 5607 4872 6983 5668
rect 11248 5035 12527 5731
rect 11246 4832 12534 5035
rect 6539 4493 9717 4590
rect 3050 4395 6089 4493
rect 3027 3791 6089 4395
rect 6538 3791 9717 4493
rect 3027 3786 5613 3791
rect 3027 3773 4434 3786
rect 7344 3763 9717 3791
rect 7344 3743 7765 3763
<< pwell >>
rect 10347 3639 13243 4492
rect 4679 2204 5969 3004
rect 6578 2204 7810 3004
<< nmos >>
rect 10469 4134 12989 4187
rect 4922 2686 5921 2742
rect 6625 2679 7624 2735
<< mvpmos >>
rect 5797 5336 6801 5391
rect 11369 5354 12385 5411
rect 3497 4134 6009 4186
rect 6629 4142 9141 4194
<< ndiff >>
rect 10469 4358 12989 4392
rect 10469 4353 12449 4358
rect 10469 4267 10535 4353
rect 10994 4348 12449 4353
rect 10994 4267 11480 4348
rect 10469 4262 11480 4267
rect 11939 4272 12449 4348
rect 12908 4272 12989 4358
rect 11939 4262 12989 4272
rect 10469 4187 12989 4262
rect 10469 4050 12989 4134
rect 10469 4040 11475 4050
rect 10469 3954 10530 4040
rect 10989 3964 11475 4040
rect 11934 3964 12449 4050
rect 12908 3964 12989 4050
rect 10989 3954 12989 3964
rect 10469 3916 12989 3954
rect 4922 2865 5921 2943
rect 4922 2814 4987 2865
rect 5209 2814 5626 2865
rect 5848 2814 5921 2865
rect 4922 2742 5921 2814
rect 6625 2858 7624 2936
rect 6625 2807 6690 2858
rect 6912 2807 7329 2858
rect 7551 2807 7624 2858
rect 6625 2735 7624 2807
rect 4922 2607 5921 2686
rect 8207 2733 8227 2734
rect 8207 2715 8208 2733
rect 8226 2715 8227 2733
rect 8207 2714 8227 2715
rect 4922 2522 4991 2607
rect 5213 2522 5607 2607
rect 5829 2522 5921 2607
rect 4922 2488 5921 2522
rect 6625 2600 7624 2679
rect 8278 2733 8297 2734
rect 8278 2715 8279 2733
rect 8296 2715 8297 2733
rect 8278 2714 8297 2715
rect 6625 2515 6694 2600
rect 6916 2515 7310 2600
rect 7532 2515 7624 2600
rect 6625 2481 7624 2515
<< mvpdiff >>
rect 5797 5685 6801 5747
rect 5797 5497 5855 5685
rect 6043 5673 6801 5685
rect 6043 5497 6575 5673
rect 5797 5485 6575 5497
rect 6763 5485 6801 5673
rect 11369 5651 12385 5731
rect 5797 5391 6801 5485
rect 11369 5532 11436 5651
rect 11760 5532 11988 5651
rect 12312 5532 12385 5651
rect 11369 5411 12385 5532
rect 5797 5269 6801 5336
rect 5797 5257 6567 5269
rect 5797 5069 5855 5257
rect 6043 5081 6567 5257
rect 6755 5081 6801 5269
rect 6043 5069 6801 5081
rect 5797 5030 6801 5069
rect 11369 5246 12385 5354
rect 11369 5231 12003 5246
rect 11369 5112 11436 5231
rect 11760 5127 12003 5231
rect 12327 5127 12385 5246
rect 11760 5112 12385 5127
rect 11369 5040 12385 5112
rect 3497 4334 6009 4392
rect 3497 4322 4433 4334
rect 3497 4237 3551 4322
rect 4079 4249 4433 4322
rect 4961 4332 6009 4334
rect 4961 4249 5426 4332
rect 4079 4247 5426 4249
rect 5954 4247 6009 4332
rect 4079 4237 6009 4247
rect 3497 4186 6009 4237
rect 6629 4342 9141 4400
rect 6629 4330 7565 4342
rect 6629 4245 6683 4330
rect 7211 4257 7565 4330
rect 8093 4340 9141 4342
rect 8093 4257 8558 4340
rect 7211 4255 8558 4257
rect 9086 4255 9141 4340
rect 7211 4245 9141 4255
rect 6629 4194 9141 4245
rect 3497 4070 6009 4134
rect 3497 4066 5430 4070
rect 3497 3981 3551 4066
rect 4079 4060 5430 4066
rect 4079 3981 4441 4060
rect 3497 3975 4441 3981
rect 4969 3985 5430 4060
rect 5958 3985 6009 4070
rect 4969 3975 6009 3985
rect 3497 3932 6009 3975
rect 6629 4078 9141 4142
rect 6629 4074 8562 4078
rect 6629 3989 6683 4074
rect 7211 4068 8562 4074
rect 7211 3989 7573 4068
rect 6629 3983 7573 3989
rect 8101 3993 8562 4068
rect 9090 3993 9141 4078
rect 8101 3983 9141 3993
rect 6629 3940 9141 3983
<< ndiffc >>
rect 10535 4267 10994 4353
rect 11480 4262 11939 4348
rect 12449 4272 12908 4358
rect 10530 3954 10989 4040
rect 11475 3964 11934 4050
rect 12449 3964 12908 4050
rect 4987 2814 5209 2865
rect 5626 2814 5848 2865
rect 6690 2807 6912 2858
rect 7329 2807 7551 2858
rect 8208 2715 8226 2733
rect 4991 2522 5213 2607
rect 5607 2522 5829 2607
rect 8279 2715 8296 2733
rect 6694 2515 6916 2600
rect 7310 2515 7532 2600
<< mvpdiffc >>
rect 5855 5497 6043 5685
rect 6575 5485 6763 5673
rect 11436 5532 11760 5651
rect 11988 5532 12312 5651
rect 5855 5069 6043 5257
rect 6567 5081 6755 5269
rect 11436 5112 11760 5231
rect 12003 5127 12327 5246
rect 3551 4237 4079 4322
rect 4433 4249 4961 4334
rect 5426 4247 5954 4332
rect 6683 4245 7211 4330
rect 7565 4257 8093 4342
rect 8558 4255 9086 4340
rect 3551 3981 4079 4066
rect 4441 3975 4969 4060
rect 5430 3985 5958 4070
rect 6683 3989 7211 4074
rect 7573 3983 8101 4068
rect 8562 3993 9090 4078
<< psubdiff >>
rect 10463 3844 12985 3889
rect 10463 3758 10525 3844
rect 10984 3758 11480 3844
rect 11939 3758 12454 3844
rect 12913 3758 12985 3844
rect 10463 3713 12985 3758
rect 4915 2398 5917 2440
rect 4915 2312 4981 2398
rect 5203 2395 5917 2398
rect 5203 2312 5609 2395
rect 4915 2309 5609 2312
rect 5831 2309 5917 2395
rect 4915 2238 5917 2309
rect 6618 2391 7620 2433
rect 6618 2305 6684 2391
rect 6906 2388 7620 2391
rect 6906 2305 7312 2388
rect 6618 2302 7312 2305
rect 7534 2302 7620 2388
rect 6618 2237 7620 2302
<< nsubdiff >>
rect 11367 5960 12385 6045
rect 11367 5812 11478 5960
rect 11673 5956 12385 5960
rect 11673 5812 12049 5956
rect 11367 5808 12049 5812
rect 12244 5808 12385 5956
rect 11367 5760 12385 5808
<< mvnsubdiff >>
rect 5797 6076 6801 6130
rect 5797 6072 6539 6076
rect 5797 5884 5867 6072
rect 6055 5888 6539 6072
rect 6727 5888 6801 6076
rect 6055 5884 6801 5888
rect 5797 5787 6801 5884
<< psubdiffcont >>
rect 10525 3758 10984 3844
rect 11480 3758 11939 3844
rect 12454 3758 12913 3844
rect 4981 2312 5203 2398
rect 5609 2309 5831 2395
rect 6684 2305 6906 2391
rect 7312 2302 7534 2388
<< nsubdiffcont >>
rect 11478 5812 11673 5960
rect 12049 5808 12244 5956
<< mvnsubdiffcont >>
rect 5867 5884 6055 6072
rect 6539 5888 6727 6076
<< poly >>
rect 9020 5566 9270 5627
rect 9020 5437 9080 5566
rect 9217 5437 9270 5566
rect 9020 5410 9270 5437
rect 11289 5411 11333 5413
rect 11289 5410 11369 5411
rect 6901 5409 11369 5410
rect 6838 5391 11369 5409
rect 5724 5336 5797 5391
rect 6801 5354 11369 5391
rect 12385 5354 12483 5411
rect 6801 5336 11329 5354
rect 6838 5332 11329 5336
rect 6838 5329 11300 5332
rect 6901 5327 11300 5329
rect 9020 5323 9270 5327
rect 3104 4249 3351 4297
rect 3104 4130 3138 4249
rect 3325 4218 3351 4249
rect 3325 4186 3446 4218
rect 9303 4281 9550 4305
rect 9303 4234 9353 4281
rect 9199 4194 9353 4234
rect 3325 4134 3497 4186
rect 6009 4134 6052 4186
rect 6578 4142 6629 4194
rect 9141 4162 9353 4194
rect 9540 4162 9550 4281
rect 9141 4142 9550 4162
rect 3325 4130 3446 4134
rect 3104 4098 3446 4130
rect 3104 4042 3351 4098
rect 9199 4114 9550 4142
rect 10079 4208 10435 4249
rect 10079 4156 10112 4208
rect 10198 4187 10435 4208
rect 10198 4156 10469 4187
rect 10079 4134 10469 4156
rect 12989 4134 13032 4187
rect 10079 4119 10435 4134
rect 10079 4115 10383 4119
rect 9303 4050 9550 4114
rect 6114 2763 6245 2783
rect 4814 2686 4922 2742
rect 5921 2736 5969 2742
rect 6114 2736 6139 2763
rect 5921 2721 6139 2736
rect 6216 2736 6245 2763
rect 6216 2735 6610 2736
rect 6216 2721 6625 2735
rect 5921 2688 6625 2721
rect 5921 2686 5969 2688
rect 6578 2679 6625 2688
rect 7624 2679 7721 2735
<< polycont >>
rect 9080 5437 9217 5566
rect 3138 4130 3325 4249
rect 9353 4162 9540 4281
rect 10112 4156 10198 4208
rect 6139 2721 6216 2763
<< ndiffres >>
rect 8197 2734 8237 2744
rect 8197 2714 8207 2734
rect 8227 2714 8237 2734
rect 8197 2673 8237 2714
rect 8266 2734 8307 2745
rect 8266 2714 8278 2734
rect 8297 2714 8307 2734
rect 8266 2705 8307 2714
rect 8267 2673 8307 2705
rect 8197 2644 8307 2673
<< locali >>
rect 5798 6127 6804 6136
rect 5798 6123 6983 6127
rect 5798 6076 11138 6123
rect 5798 6072 6539 6076
rect 5798 5884 5867 6072
rect 6055 6065 6539 6072
rect 6727 6065 11138 6076
rect 6055 5903 6532 6065
rect 6730 6045 11138 6065
rect 11367 6045 12385 6049
rect 6730 5960 12385 6045
rect 6730 5903 11478 5960
rect 6055 5888 6539 5903
rect 6727 5888 11478 5903
rect 6055 5884 11478 5888
rect 5798 5883 11138 5884
rect 5798 5881 6983 5883
rect 5798 5685 6804 5881
rect 5798 5674 5855 5685
rect 6043 5674 6804 5685
rect 5798 5512 5848 5674
rect 6046 5673 6804 5674
rect 6046 5658 6575 5673
rect 6763 5658 6804 5673
rect 6046 5512 6572 5658
rect 5798 5497 5855 5512
rect 6043 5497 6572 5512
rect 5798 5496 6572 5497
rect 6770 5496 6804 5658
rect 11365 5812 11478 5884
rect 11673 5956 12385 5960
rect 11673 5812 12049 5956
rect 11365 5808 12049 5812
rect 12244 5808 12385 5956
rect 11365 5753 12385 5808
rect 11365 5654 12388 5753
rect 11365 5651 11440 5654
rect 5798 5485 6575 5496
rect 6763 5485 6804 5496
rect 5798 5417 6804 5485
rect 9020 5566 9270 5627
rect 9020 5437 9080 5566
rect 9217 5437 9270 5566
rect 11365 5532 11436 5651
rect 11365 5531 11440 5532
rect 11760 5531 11987 5654
rect 12310 5651 12388 5654
rect 12312 5532 12388 5651
rect 12310 5531 12388 5532
rect 11365 5458 12388 5531
rect 9020 5323 9270 5437
rect 5798 5269 6800 5309
rect 5798 5257 6567 5269
rect 5798 5069 5855 5257
rect 6043 5081 6567 5257
rect 6755 5081 6800 5269
rect 6043 5069 6800 5081
rect 5798 5053 6800 5069
rect 11370 5257 12394 5316
rect 11370 5246 12399 5257
rect 11370 5231 12003 5246
rect 11370 5112 11436 5231
rect 11760 5127 12003 5231
rect 12327 5127 12399 5246
rect 11760 5112 12399 5127
rect 5782 5021 6856 5053
rect 11370 5042 12399 5112
rect 5782 4933 6009 5021
rect 5740 4493 6009 4933
rect 6629 4941 6856 5021
rect 6629 4872 6904 4941
rect 6635 4493 6904 4872
rect 12111 4816 12399 5042
rect 12111 4815 13176 4816
rect 13388 4815 13505 4820
rect 12111 4627 13505 4815
rect 5717 4442 6009 4493
rect 5717 4397 6004 4442
rect 3507 4353 6004 4397
rect 6633 4405 6920 4493
rect 6633 4353 9134 4405
rect 12444 4398 12732 4627
rect 13150 4624 13505 4627
rect 3507 4334 6002 4353
rect 3507 4322 4433 4334
rect 3096 4249 3367 4297
rect 3096 4130 3138 4249
rect 3325 4130 3367 4249
rect 3507 4237 3551 4322
rect 4079 4249 4433 4322
rect 4961 4332 6002 4334
rect 4961 4249 5426 4332
rect 4079 4247 5426 4249
rect 5954 4247 6002 4332
rect 4079 4237 6002 4247
rect 3507 4206 6002 4237
rect 6639 4342 9134 4353
rect 6639 4330 7565 4342
rect 6639 4245 6683 4330
rect 7211 4257 7565 4330
rect 8093 4340 9134 4342
rect 8093 4257 8558 4340
rect 7211 4255 8558 4257
rect 9086 4255 9134 4340
rect 10473 4358 12990 4398
rect 10473 4353 12449 4358
rect 7211 4245 9134 4255
rect 6639 4214 9134 4245
rect 9287 4281 9558 4305
rect 3096 4042 3367 4130
rect 9287 4162 9353 4281
rect 9540 4162 9558 4281
rect 10473 4267 10535 4353
rect 10994 4348 12449 4353
rect 10994 4267 11480 4348
rect 10473 4262 11480 4267
rect 11939 4272 12449 4348
rect 12908 4272 12990 4358
rect 11939 4262 12990 4272
rect 3511 4070 6006 4119
rect 3511 4066 5430 4070
rect 3511 3981 3551 4066
rect 4079 4060 5430 4066
rect 4079 3981 4441 4060
rect 3511 3975 4441 3981
rect 4969 3985 5430 4060
rect 5958 3985 6006 4070
rect 4969 3975 6006 3985
rect 3511 3928 6006 3975
rect 6643 4078 9138 4127
rect 6643 4074 8562 4078
rect 6643 3989 6683 4074
rect 7211 4068 8562 4074
rect 7211 3989 7573 4068
rect 6643 3983 7573 3989
rect 8101 3993 8562 4068
rect 9090 3993 9138 4078
rect 9287 4050 9558 4162
rect 10079 4208 10235 4254
rect 10473 4227 12990 4262
rect 13388 4233 13505 4624
rect 10079 4156 10112 4208
rect 10198 4156 10235 4208
rect 8101 3983 9138 3993
rect 6643 3936 9138 3983
rect 5757 3840 5916 3928
rect 5747 3791 5916 3840
rect 6713 3829 6857 3936
rect 6708 3811 6861 3829
rect 6708 3791 6869 3811
rect 5747 3213 5915 3791
rect 6708 3417 6861 3791
rect 8191 3632 8238 3637
rect 10079 3632 10235 4156
rect 13388 4166 13412 4233
rect 13479 4166 13505 4233
rect 10463 4050 12985 4095
rect 10463 4040 11475 4050
rect 10463 3954 10530 4040
rect 10989 3964 11475 4040
rect 11934 3964 12449 4050
rect 12908 3964 12985 4050
rect 10989 3954 12985 3964
rect 10463 3848 12985 3954
rect 10463 3844 10532 3848
rect 10981 3845 12985 3848
rect 10981 3844 11481 3845
rect 11931 3844 12463 3845
rect 10463 3758 10525 3844
rect 10984 3758 11480 3844
rect 11939 3758 12454 3844
rect 10463 3756 11481 3758
rect 11931 3756 12463 3758
rect 12913 3756 12985 3845
rect 10463 3713 12985 3756
rect 8191 3559 10239 3632
rect 6707 3416 7597 3417
rect 8191 3416 8238 3559
rect 12139 3459 12351 3460
rect 13388 3459 13505 4166
rect 11295 3427 11759 3430
rect 11244 3424 11759 3427
rect 6707 3277 8239 3416
rect 9875 3395 11759 3424
rect 9875 3374 11477 3395
rect 11498 3374 11759 3395
rect 9875 3351 11759 3374
rect 12139 3429 13505 3459
rect 12139 3411 12165 3429
rect 12182 3411 12201 3429
rect 12218 3411 12237 3429
rect 12254 3411 12273 3429
rect 12290 3411 13505 3429
rect 12139 3379 13505 3411
rect 12139 3373 12371 3379
rect 12139 3370 12351 3373
rect 6707 3267 7597 3277
rect 6708 3220 6861 3267
rect 5747 3182 5919 3213
rect 6708 3201 6869 3220
rect 5749 3166 5919 3182
rect 5749 3163 6238 3166
rect 5749 3057 6245 3163
rect 5749 2910 5903 3057
rect 4952 2888 5903 2910
rect 4952 2865 5894 2888
rect 4952 2814 4987 2865
rect 5209 2814 5626 2865
rect 5848 2814 5894 2865
rect 4952 2776 5894 2814
rect 6114 2763 6245 3057
rect 6715 2903 6869 3201
rect 6655 2858 7597 2903
rect 6655 2807 6690 2858
rect 6912 2807 7329 2858
rect 7551 2807 7597 2858
rect 6655 2769 7597 2807
rect 6114 2721 6139 2763
rect 6216 2721 6245 2763
rect 8196 2733 8238 3277
rect 9885 3257 9922 3351
rect 11244 3347 11759 3351
rect 11295 3345 11759 3347
rect 9890 2747 9917 3257
rect 8313 2746 9922 2747
rect 8196 2724 8208 2733
rect 6114 2686 6245 2721
rect 8197 2715 8208 2724
rect 8226 2724 8238 2733
rect 8267 2733 9922 2746
rect 8226 2715 8237 2724
rect 8197 2704 8237 2715
rect 8267 2715 8279 2733
rect 8296 2715 9922 2733
rect 8267 2711 9922 2715
rect 8267 2706 8330 2711
rect 8267 2705 8329 2706
rect 11116 2674 11213 2784
rect 4941 2607 5894 2660
rect 4941 2522 4991 2607
rect 5213 2522 5607 2607
rect 5829 2522 5894 2607
rect 4941 2398 5894 2522
rect 4941 2312 4981 2398
rect 5203 2396 5894 2398
rect 5203 2395 5620 2396
rect 5818 2395 5894 2396
rect 5203 2312 5609 2395
rect 4941 2307 4994 2312
rect 5191 2309 5609 2312
rect 5831 2309 5894 2395
rect 5191 2307 5620 2309
rect 5818 2307 5894 2309
rect 4941 2260 5894 2307
rect 6644 2600 7597 2653
rect 6644 2515 6694 2600
rect 6916 2515 7310 2600
rect 7532 2515 7597 2600
rect 6644 2393 7597 2515
rect 6644 2391 6701 2393
rect 6898 2391 7322 2393
rect 6644 2305 6684 2391
rect 6906 2388 7322 2391
rect 7519 2388 7597 2393
rect 6906 2305 7312 2388
rect 6644 2303 6701 2305
rect 6898 2303 7312 2305
rect 6644 2302 7312 2303
rect 7534 2302 7597 2388
rect 6644 2253 7597 2302
<< viali >>
rect 5878 5897 6040 6059
rect 6532 5903 6539 6065
rect 6539 5903 6727 6065
rect 6727 5903 6730 6065
rect 5848 5512 5855 5674
rect 5855 5512 6043 5674
rect 6043 5512 6046 5674
rect 6572 5496 6575 5658
rect 6575 5496 6763 5658
rect 6763 5496 6770 5658
rect 11478 5812 11673 5960
rect 12049 5808 12244 5956
rect 11440 5651 11760 5654
rect 11440 5532 11760 5651
rect 11440 5531 11760 5532
rect 11987 5651 12310 5654
rect 11987 5532 11988 5651
rect 11988 5532 12310 5651
rect 11987 5531 12310 5532
rect 13412 4166 13479 4233
rect 10532 3844 10981 3848
rect 11481 3844 11931 3845
rect 12463 3844 12913 3845
rect 10532 3758 10981 3844
rect 11481 3758 11931 3844
rect 12463 3758 12913 3844
rect 11481 3756 11931 3758
rect 12463 3756 12913 3758
rect 11477 3374 11498 3395
rect 12165 3411 12182 3429
rect 12201 3411 12218 3429
rect 12237 3411 12254 3429
rect 12273 3411 12290 3429
rect 4994 2312 5191 2396
rect 5620 2395 5818 2396
rect 4994 2307 5191 2312
rect 5620 2309 5818 2395
rect 5620 2307 5818 2309
rect 6701 2391 6898 2393
rect 6701 2305 6898 2391
rect 7322 2388 7519 2393
rect 6701 2303 6898 2305
rect 7322 2303 7519 2388
<< metal1 >>
rect 6166 6120 6418 6749
rect 5758 6065 6832 6120
rect 5758 6059 6532 6065
rect 5758 5897 5878 6059
rect 6040 5903 6532 6059
rect 6730 5903 6832 6065
rect 6040 5897 6832 5903
rect 5758 5674 6832 5897
rect 5758 5512 5848 5674
rect 6046 5658 6832 5674
rect 6046 5512 6572 5658
rect 5758 5496 6572 5512
rect 6770 5496 6832 5658
rect 5758 5445 6832 5496
rect 9677 4913 9914 6675
rect 11360 5960 12388 6048
rect 11360 5812 11478 5960
rect 11673 5956 12388 5960
rect 11673 5812 12049 5956
rect 11360 5808 12049 5812
rect 12244 5808 12388 5956
rect 11360 5654 12388 5808
rect 11360 5531 11440 5654
rect 11760 5531 11987 5654
rect 12310 5531 12388 5654
rect 11360 5458 12388 5531
rect 9306 4691 9914 4913
rect 2538 4009 3353 4291
rect 9306 4039 9558 4691
rect 13386 4233 13676 4267
rect 13386 4166 13412 4233
rect 13479 4166 13676 4233
rect 13386 4140 13676 4166
rect 10429 3874 13019 4085
rect 7877 3848 13019 3874
rect 7877 3758 10532 3848
rect 10981 3845 13019 3848
rect 10981 3758 11481 3845
rect 7877 3756 11481 3758
rect 11931 3756 12463 3845
rect 12913 3756 13019 3845
rect 7877 3732 13019 3756
rect 7877 3692 10530 3732
rect 4861 2640 5969 2647
rect 4852 2526 5969 2640
rect 6578 2526 7675 2640
rect 4852 2413 7675 2526
rect 7885 2413 7998 3692
rect 10323 2784 10371 3692
rect 11303 3395 11762 3430
rect 11303 3374 11477 3395
rect 11498 3374 11762 3395
rect 11303 3345 11762 3374
rect 12139 3429 12316 3463
rect 12139 3411 12165 3429
rect 12182 3411 12201 3429
rect 12218 3411 12237 3429
rect 12254 3411 12273 3429
rect 12290 3411 12316 3429
rect 12139 3370 12316 3411
rect 10321 2781 11069 2784
rect 10321 2779 11074 2781
rect 10321 2737 11206 2779
rect 10321 2711 11151 2737
rect 11178 2711 11206 2737
rect 10321 2678 11206 2711
rect 10323 2654 10371 2678
rect 11037 2677 11206 2678
rect 4852 2402 7998 2413
rect 4852 2396 5969 2402
rect 4852 2307 4994 2396
rect 5191 2307 5620 2396
rect 5818 2307 5969 2396
rect 4852 2269 5969 2307
rect 4861 2263 5969 2269
rect 6578 2393 7998 2402
rect 6578 2303 6701 2393
rect 6898 2303 7322 2393
rect 7519 2303 7998 2393
rect 6578 2258 7998 2303
rect 6578 2256 7675 2258
rect 7874 1779 7994 2258
<< via1 >>
rect 11151 2711 11178 2737
<< metal2 >>
rect 12286 3313 12311 3320
rect 11309 3310 11763 3313
rect 12001 3310 12311 3313
rect 11214 3303 12311 3310
rect 11214 3302 12309 3303
rect 11214 2781 12307 3302
rect 11114 2737 12307 2781
rect 11114 2711 11151 2737
rect 11178 2711 12307 2737
rect 11114 2677 12307 2711
rect 11214 2222 12307 2677
<< metal3 >>
rect 12141 3313 12309 3458
rect 12001 3310 12311 3313
rect 11214 2957 12311 3310
rect 11214 2222 12307 2957
<< mimcap >>
rect 11260 3162 12259 3267
rect 11260 2810 11353 3162
rect 11705 3161 12259 3162
rect 11708 2811 12259 3161
rect 11705 2810 12259 2811
rect 11260 2268 12259 2810
<< mimcapcontact >>
rect 11353 3161 11705 3162
rect 11353 2811 11708 3161
rect 11353 2810 11705 2811
<< metal4 >>
rect 11308 3313 11759 3428
rect 11308 3298 11763 3313
rect 11310 3162 11763 3298
rect 11310 2810 11353 3162
rect 11705 3161 11763 3162
rect 11708 2811 11763 3161
rect 11705 2810 11763 2811
rect 11310 2742 11763 2810
use pmos_substrate  pmos_substrate_3
timestamp 1633808399
transform 1 0 11825 0 1 4928
box -33 -34 81 81
use pmos_substrate  pmos_substrate_2
timestamp 1633808399
transform 1 0 7860 0 1 4483
box -33 -34 81 81
use pmos_substrate  pmos_substrate_1
timestamp 1633808399
transform 1 0 4736 0 1 3827
box -33 -34 81 81
use pmos_substrate  pmos_substrate_0
timestamp 1633808399
transform 1 0 6291 0 1 4928
box -33 -34 81 81
use nmos_substrate  nmos_substrate_2
timestamp 1633808399
transform 1 0 7681 0 1 2900
box 0 0 48 48
use nmos_substrate  nmos_substrate_1
timestamp 1633808399
transform 1 0 4765 0 1 2831
box 0 0 48 48
use nmos_substrate  nmos_substrate_0
timestamp 1633808399
transform 1 0 13111 0 1 3787
box 0 0 48 48
<< labels >>
rlabel metal1 s 5236 2276 5292 2414 4 gnd
rlabel locali s 6771 3074 6821 3206 4 vo
rlabel locali s 3136 4042 3311 4098 4 vinp
rlabel locali s 9358 4058 9533 4114 4 vinm
rlabel metal1 s 5876 5787 6053 5851 4 vdd
rlabel locali s 13397 4071 13491 4116 4 vout
rlabel locali s 10234 3371 10304 3401 4 top
rlabel metal4 s 11452 3351 11525 3364 4 top
rlabel metal3 s 12192 3379 12249 3394 4 vout
rlabel metal2 s 11136 2761 11181 2779 4 gnd
rlabel locali 9073 5346 9202 5392 1 vbias
rlabel locali 6152 2692 6199 2709 1 vg
<< properties >>
string FIXED_BBOX 0 0 5672 4169
<< end >>
